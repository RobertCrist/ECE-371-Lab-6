module playerControl();

endmodule
